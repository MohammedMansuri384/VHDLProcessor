library verilog;
use verilog.vl_types.all;
entity ModALU_vlg_vec_tst is
end ModALU_vlg_vec_tst;
